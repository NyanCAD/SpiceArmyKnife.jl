Diode cascade (Voltage multiplier)

vs a 0 dc=0 sin 0 50 100k
r1 a 1 0.01
c1 1 2 100n
xd1 0 1 sp_diode is=76.9p rs=42.0m cjo=26.5p m=0.333 n=1.45 tt=4.32u
c2 0 10 100n
xd2 1 10 sp_diode is=76.9p rs=42.0m cjo=26.5p m=0.333 n=1.45 tt=4.32u
c3 1 2 100n
xd3 10 2 sp_diode is=76.9p rs=42.0m cjo=26.5p m=0.333 n=1.45 tt=4.32u
c4 10 20 100n
xd4 2 20 sp_diode is=76.9p rs=42.0m cjo=26.5p m=0.333 n=1.45 tt=4.32u

.end
