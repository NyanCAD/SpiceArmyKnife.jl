RC circuit excited by a pulse train

vs 1 0 dc 0 pulse 0 1 1u 1u 1u 1m 2m
r1 1 2 1k
c1 2 0 1u

.tran 1u 1 0 1u

.end
